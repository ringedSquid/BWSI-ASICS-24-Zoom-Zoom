`default_nettype none

module alu (

);

endmodule
